module AND (Entrada1, Entrada2, Resultado);

  input Entrada1, Entrada2;
  output Resultado;

  assign Resultado = Entrada1 & Entrada2;

endmodule
